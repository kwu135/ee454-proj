module tb_HuffmanEncode();

reg clk, start, reset;
reg [95:0] data_in0;
reg [95:0] data_in1;
reg [95:0] data_in2;
reg [95:0] data_in3;
reg [95:0] data_in4;
reg [95:0] data_in5;
reg [95:0] data_in6;
reg [95:0] data_in7;

wire [8:0] num_bits;
wire done;
wire [511:0] data_out;
parameter CLK_PERIOD=2;
always 	#(CLK_PERIOD/2) clk=~clk;

initial 
begin
clk=0;
reset =0;
/*
data_in0 = 
12'b111111111101 << 84 |
12'b000000000000 << 72 |
12'b111111110101 << 60 |
12'b000000001001 << 48 |
12'b000000000101 << 36 |
12'b000000000111 << 24 |
12'b111111111000 << 12 |
12'b000000000100;

data_in1 = 
12'b000000000001<< 84 |
12'b000000000100 << 72 |
12'b000000000000 << 60 |
12'b111111111111 << 48 |
12'b000000000001 << 36 |
12'b111111110101 << 24 |
12'b000000000011 << 12 |
12'b111111010001;

data_in2 = 
12'b000000000110<< 84 |
12'b000000000100<< 72 |
12'b111111111101<< 60 |
12'b000000000001 << 48 |
12'b000000000101 << 36 |
12'b111111110100 << 24 |
12'b000000001001 << 12 |
12'b000000000101;
data_in3 = 
12'b000000000001<< 84 |
12'b000000000100 << 72 |
12'b000000000000 << 60 |
12'b111111111111 << 48 |
12'b000000000001 << 36 |
12'b111111110101 << 24 |
12'b000000000011 << 12 |
12'b111111010001;
data_in4 = 
12'b000000000001<< 84 |
12'b000000000100 << 72 |
12'b000000000000 << 60 |
12'b111111111111 << 48 |
12'b000000000001 << 36 |
12'b111111110101 << 24 |
12'b000000000011 << 12 |
12'b111111010001;
data_in5 = 
12'b000000000001<< 84 |
12'b000000000100 << 72 |
12'b000000000000 << 60 |
12'b111111111111 << 48 |
12'b000000000001 << 36 |
12'b111111110101 << 24 |
12'b000000000011 << 12 |
12'b111111010001;
data_in6 = 
12'b000000000001<< 84 |
12'b000000000100 << 72 |
12'b000000000000 << 60 |
12'b111111111111 << 48 |
12'b000000000001 << 36 |
12'b111111110101 << 24 |
12'b000000000011 << 12 |
12'b111111010001;
data_in7 = 
12'b000000000001<< 84 |
12'b000000000100 << 72 |
12'b000000000000 << 60 |
12'b111111111111 << 48 |
12'b000000000001 << 36 |
12'b111111110101 << 24 |
12'b000000000011 << 12 |
12'b111111010001; */

data_in0 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000100;

data_in1 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;

data_in2 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;
data_in3 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;
data_in4 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;
data_in5 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;
data_in6 = 
12'b000000000000 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;
data_in7 = 
12'b111111111111 << 84 |
12'b000000000000 << 72 |
12'b000000000000 << 60 |
12'b000000000000 << 48 |
12'b000000000000 << 36 |
12'b000000000000 << 24 |
12'b000000000000 << 12 |
12'b000000000000;


#(CLK_PERIOD*5)
reset = 1;
#(CLK_PERIOD)
reset = 0;
#(CLK_PERIOD)
start = 1;
#(CLK_PERIOD * 80)
$stop;
end

HuffmanEncode encoder(clk, data_in0, data_in1, data_in2, data_in3, data_in4,
	data_in5, data_in6, data_in7, reset, start, data_out, num_bits, done);
endmodule // tb_HuffmanEncode
