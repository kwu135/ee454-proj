module Quant(in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, clk, 
	q_0,q_1,q_2,q_3,q_4,q_5,q_6,q_7);
  
input [95:0] in_0; 
input [95:0] in_1; 
input [95:0] in_2; 
input [95:0] in_3; 
input [95:0] in_4; 
input [95:0] in_5; 
input [95:0] in_6; 
input [95:0] in_7; 
input clk;
output [95:0] q_0; reg [95:0]q_0;
output [95:0] q_1; reg [95:0]q_1;
output [95:0] q_2; reg [95:0]q_2;
output [95:0] q_3; reg [95:0]q_3;
output [95:0] q_4; reg [95:0]q_4;
output [95:0] q_5; reg [95:0]q_5;
output [95:0] q_6; reg [95:0]q_6;
output [95:0] q_7; reg [95:0]q_7;
reg [7:0] Quant [7:0][7:0];


	initial begin
	Quant[0][0]<= 16;
	Quant[0][1]<= 11;
	Quant[0][2]<= 10;
	Quant[0][3]<= 16;
	Quant[0][4]<= 24;
	Quant[0][5]<= 40;
	Quant[0][6]<= 51;
	Quant[0][7]<= 61;
	Quant[1][0]<= 12;
	Quant[1][1]<= 12;
	Quant[1][2]<= 14;
	Quant[1][3]<= 19;
	Quant[1][4]<= 26;
	Quant[1][5]<= 58;
	Quant[1][6]<= 60;
	Quant[1][7]<= 55;
	Quant[2][0]<= 14;
	Quant[2][1]<= 13;
	Quant[2][2]<= 16;
	Quant[2][3]<= 24;
	Quant[2][4]<= 40;
	Quant[2][5]<= 57;
	Quant[2][6]<= 69;
	Quant[2][7]<= 56;
	Quant[3][0]<= 14;
	Quant[3][1]<= 17;
	Quant[3][2]<= 22;
	Quant[3][3]<= 29;
	Quant[3][4]<= 51;
	Quant[3][5]<= 87;
	Quant[3][6]<= 80;
	Quant[3][7]<= 62;
	Quant[4][0]<= 18;
	Quant[4][1]<= 22;
	Quant[4][2]<= 37;
	Quant[4][3]<= 56;
	Quant[4][4]<= 68;
	Quant[4][5]<= 109;
	Quant[4][6]<= 103;
	Quant[4][7]<= 77;
	Quant[5][0]<= 24;
	Quant[5][1]<= 35;
	Quant[5][2]<= 55;
	Quant[5][3]<= 64;
	Quant[5][4]<= 81;
	Quant[5][5]<= 104;
	Quant[5][6]<= 113;
	Quant[5][7]<= 92;
	Quant[6][0]<= 49;
	Quant[6][1]<= 64;
	Quant[6][2]<= 78;
	Quant[6][3]<= 87;
	Quant[6][4]<= 103;
	Quant[6][5]<= 121;
	Quant[6][6]<= 120;
	Quant[6][7]<= 101;
	Quant[7][0]<= 72;
	Quant[7][1]<= 92;
	Quant[7][2]<= 95;
	Quant[7][3]<= 98;
	Quant[7][4]<= 112;
	Quant[7][5]<= 100;
	Quant[7][6]<= 103;
	Quant[7][7]<= 99;
	end
	
	always @(posedge clk)
	begin

    	if(in_0[95:84] > 12'b011111111111)
		begin
			q_0[95:84] = ((in_0[95:84]^12'b111111111111)+1) / Quant[0][7];
			if (q_0[95:84] >0) q_0[95:84] =(q_0[95:84]^12'b111111111111)+1;
		end
		else q_0[95:84] = in_0[95:84] / Quant[0][7];

		if(in_0[83:72] > 12'b011111111111)
		begin
			q_0[83:72] = ((in_0[83:72]^12'b111111111111)+1) / Quant[0][6];
			if (q_0[83:72] >0) q_0[83:72] =(q_0[83:72]^12'b111111111111)+1;
		end
		else q_0[83:72] = in_0[83:72] / Quant[0][6];

		if(in_0[71:60] > 12'b011111111111)
		begin
			q_0[71:60] = ((in_0[71:60]^12'b111111111111)+1) / Quant[0][5];
			if (q_0[71:60] >0) q_0[71:60] =(q_0[71:60]^12'b111111111111)+1;
		end
		else q_0[71:60] = in_0[71:60] / Quant[0][5];

		if(in_0[59:48] > 12'b011111111111)
		begin
			q_0[59:48] = ((in_0[59:48]^12'b111111111111)+1) / Quant[0][4];
			if (q_0[59:48] >0) q_0[59:48] =(q_0[59:48]^12'b111111111111)+1;
		end
		else q_0[59:48] = in_0[59:48] / Quant[0][4];

		if(in_0[47:36] > 12'b011111111111)
		begin
			q_0[47:36] = ((in_0[47:36]^12'b111111111111)+1) / Quant[0][3];
			if (q_0[47:36] >0) q_0[47:36] =(q_0[47:36]^12'b111111111111)+1;
		end
		else q_0[47:36] = in_0[47:36] / Quant[0][3];

		if(in_0[35:24] > 12'b011111111111)
		begin
			q_0[35:24] = ((in_0[35:24]^12'b111111111111)+1) / Quant[0][2];
			if (q_0[35:24] >0) q_0[35:24] =(q_0[35:24]^12'b111111111111)+1;
		end
		else q_0[35:24] = in_0[35:24] / Quant[0][2];

		if(in_0[23:12] > 12'b011111111111)
		begin
			q_0[23:12] = ((in_0[23:12]^12'b111111111111)+1) / Quant[0][1];
			if (q_0[23:12] >0) q_0[23:12] =(q_0[23:12]^12'b111111111111)+1;
		end
		else q_0[23:12] = in_0[23:12] / Quant[0][1];

		if(in_0[11:0]  > 12'b011111111111)
		begin
			q_0[11:0] = ((in_0[11:0]^12'b111111111111)+1) / Quant[0][0];
			if (q_0[11:0] >0) q_0[11:0]  =(q_0[11:0])^12'b1111111111111+1;
		end
		else q_0[11:0]  = in_0[11:0] /  Quant[0][0];

		if(in_1[95:84] > 12'b011111111111)
		begin
			q_1[95:84] = ((in_1[95:84]^12'b111111111111)+1) / Quant[1][7];
			if (q_1[95:84] >0) q_1[95:84] =(q_1[95:84]^12'b111111111111)+1;
		end
		else q_1[95:84] = in_1[95:84] / Quant[1][7];
		if(in_1[83:72] > 12'b011111111111)
		begin
			q_1[83:72] = ((in_1[83:72]^12'b111111111111)+1) / Quant[1][6];
			if (q_1[83:72] >0) q_1[83:72] =(q_1[83:72]^12'b111111111111)+1;
		end
		else q_1[83:72] = in_1[83:72] / Quant[1][6];
		if(in_1[71:60] > 12'b011111111111)
		begin
			q_1[71:60] = ((in_1[71:60]^12'b111111111111)+1) / Quant[1][5];
			if (q_1[71:60] >0) q_1[71:60] =(q_1[71:60]^12'b111111111111)+1;
		end
		else q_1[71:60] = in_1[71:60] / Quant[1][5];
		if(in_1[59:48] > 12'b011111111111)
		begin
			q_1[59:48] = ((in_1[59:48]^12'b111111111111)+1) / Quant[1][4];
			if (q_1[59:48] >0) q_1[59:48] =(q_1[59:48]^12'b111111111111)+1;
		end
		else q_1[59:48] = in_1[59:48] / Quant[1][4];
		if(in_1[47:36] > 12'b011111111111)
		begin
			q_1[47:36] = ((in_1[47:36]^12'b111111111111)+1) / Quant[1][3];
			if (q_1[47:36] >0) q_1[47:36] =(q_1[47:36]^12'b111111111111)+1;
		end
		else q_1[47:36] = in_1[47:36] / Quant[1][3];
		if(in_1[35:24] > 12'b011111111111)
		begin
			q_1[35:24] = ((in_1[35:24]^12'b111111111111)+1) / Quant[1][2];
			if (q_1[35:24] >0) q_1[35:24] =(q_1[35:24]^12'b111111111111)+1;
		end
		else q_1[35:24] = in_1[35:24] / Quant[1][2];
		if(in_1[23:12] > 12'b011111111111)
		begin
			q_1[23:12] = ((in_1[23:12]^12'b111111111111)+1) / Quant[1][1];
			if (q_1[23:12] >0) q_1[23:12] =(q_1[23:12]^12'b111111111111)+1;
		end
		else q_1[23:12] = in_1[23:12] / Quant[1][1];
		if(in_1[11:0]  > 12'b011111111111)
		begin
			q_1[11:0]  = ((in_1[11:0] ^12'b111111111111)+1) / Quant[1][0];
			if (q_1[11:0]  >0) q_1[11:0]  =(q_1[11:0] ^12'b111111111111)+1;
		end
		else q_1[11:0]  = in_1[11:0]  / Quant[1][0];
		

		if(in_2[95:84] > 12'b011111111111)
		begin
			q_2[95:84] = ((in_2[95:84]^12'b111111111111)+1) / Quant[2][7];
			if (q_2[95:84] >0) q_2[95:84] =(q_2[95:84]^12'b111111111111)+1;
		end
		else q_2[95:84] = in_2[95:84] / Quant[2][7];
		if(in_2[83:72] > 12'b011111111111)
		begin
			q_2[83:72] = ((in_2[83:72]^12'b111111111111)+1) / Quant[2][6];
			if (q_2[83:72] >0) q_2[83:72] =(q_2[83:72]^12'b111111111111)+1;
		end
		else q_2[83:72] = in_2[83:72] / Quant[2][6];
		if(in_2[71:60] > 12'b011111111111)
		begin
			q_2[71:60] = ((in_2[71:60]^12'b111111111111)+1) / Quant[2][5];
			if (q_2[71:60] >0) q_2[71:60] =(q_2[71:60]^12'b111111111111)+1;
		end
		else q_2[71:60] = in_2[71:60] / Quant[2][5];
		if(in_2[59:48] > 12'b011111111111)
		begin
			q_2[59:48] = ((in_2[59:48]^12'b111111111111)+1) / Quant[2][4];
			if (q_2[59:48] >0) q_2[59:48] =(q_2[59:48]^12'b111111111111)+1;
		end
		else q_2[59:48] = in_2[59:48] / Quant[2][4];
		if(in_2[47:36] > 12'b011111111111)
		begin
			q_2[47:36] = ((in_2[47:36]^12'b111111111111)+1) / Quant[2][3];
			if (q_2[47:36] >0) q_2[47:36] =(q_2[47:36]^12'b111111111111)+1;
		end
		else q_2[47:36] = in_2[47:36] / Quant[2][3];
		if(in_2[35:24] > 12'b011111111111)
		begin
			q_2[35:24] = ((in_2[35:24]^12'b111111111111)+1) / Quant[2][2];
			if (q_2[35:24] >0) q_2[35:24] =(q_2[35:24]^12'b111111111111)+1;
		end
		else q_2[35:24] = in_2[35:24] / Quant[2][2];
		if(in_2[23:12] > 12'b011111111111)
		begin
			q_2[23:12] = ((in_2[23:12]^12'b111111111111)+1) / Quant[2][1];
			if (q_2[23:12] >0) q_2[23:12] =(q_2[23:12]^12'b111111111111)+1;
		end
		else q_2[23:12] = in_2[23:12] / Quant[2][1];
		if(in_2[11:0]  > 12'b011111111111)
		begin
			q_2[11:0]  = ((in_2[11:0] ^12'b111111111111)+1) / Quant[2][0];
			if (q_2[11:0]  >0) q_2[11:0]  =(q_2[11:0] ^12'b111111111111)+1;
		end
		else q_2[11:0]  = in_2[11:0]  / Quant[2][0];
		
		if(in_3[95:84] > 12'b011111111111)
		begin
			q_3[95:84] = ((in_3[95:84]^12'b111111111111)+1) / Quant[3][7];
			if (q_3[95:84] >0) q_3[95:84] =(q_3[95:84]^12'b111111111111)+1;
		end
		else q_3[95:84] = in_3[95:84] / Quant[3][7];
		if(in_3[83:72] > 12'b011111111111)
		begin
			q_3[83:72] = ((in_3[83:72]^12'b111111111111)+1) / Quant[3][6];
			if (q_3[83:72] >0) q_3[83:72] =(q_3[83:72]^12'b111111111111)+1;
		end
		else q_3[83:72] = in_3[83:72] / Quant[3][6];
		if(in_3[71:60] > 12'b011111111111)
		begin
			q_3[71:60] = ((in_3[71:60]^12'b111111111111)+1) / Quant[3][5];
			if (q_3[71:60] >0) q_3[71:60] =(q_3[71:60]^12'b111111111111)+1;
		end
		else q_3[71:60] = in_3[71:60] / Quant[3][5];
		if(in_3[59:48] > 12'b011111111111)
		begin
			q_3[59:48] = ((in_3[59:48]^12'b111111111111)+1) / Quant[3][4];
			if (q_3[59:48] >0) q_3[59:48] =(q_3[59:48]^12'b111111111111)+1;
		end
		else q_3[59:48] = in_3[59:48] / Quant[3][4];
		if(in_3[47:36] > 12'b011111111111)
		begin
			q_3[47:36] = ((in_3[47:36]^12'b111111111111)+1) / Quant[3][3];
			if (q_3[47:36] >0) q_3[47:36] =(q_3[47:36]^12'b111111111111)+1;
		end
		else q_3[47:36] = in_3[47:36] / Quant[3][3];
		if(in_3[35:24] > 12'b011111111111)
		begin
			q_3[35:24] = ((in_3[35:24]^12'b111111111111)+1) / Quant[3][2];
			if (q_3[35:24] >0) q_3[35:24] =(q_3[35:24]^12'b111111111111)+1;
		end
		else q_3[35:24] = in_3[35:24] / Quant[3][2];
		if(in_3[23:12] > 12'b011111111111)
		begin
			q_3[23:12] = ((in_3[23:12]^12'b111111111111)+1) / Quant[3][1];
			if (q_3[23:12] >0) q_3[23:12] =(q_3[23:12]^12'b111111111111)+1;
		end
		else q_3[23:12] = in_3[23:12] / Quant[3][1];
		if(in_3[11:0]  > 12'b011111111111)
		begin
			q_3[11:0]  = ((in_3[11:0] ^12'b111111111111)+1) / Quant[3][0];
			if (q_3[11:0]  >0) q_3[11:0]  =(q_3[11:0] ^12'b111111111111)+1;
		end
		else q_3[11:0]  = in_3[11:0]  / Quant[3][0];
		
		if(in_4[95:84] > 12'b011111111111)
		begin
			q_4[95:84] = ((in_4[95:84]^12'b111111111111)+1) / Quant[4][7];
			if (q_4[95:84] >0) q_4[95:84] =(q_4[95:84]^12'b111111111111)+1;
		end
		else q_4[95:84] = in_4[95:84] / Quant[4][7];
		if(in_4[83:72] > 12'b011111111111)
		begin
			q_4[83:72] = ((in_4[83:72]^12'b111111111111)+1) / Quant[4][6];
			if (q_4[83:72] >0) q_4[83:72] =(q_4[83:72]^12'b111111111111)+1;
		end
		else q_4[83:72] = in_4[83:72] / Quant[4][6];
		if(in_4[71:60] > 12'b011111111111)
		begin
			q_4[71:60] = ((in_4[71:60]^12'b111111111111)+1) / Quant[4][5];
			if (q_4[71:60] >0) q_4[71:60] =(q_4[71:60]^12'b111111111111)+1;
		end
		else q_4[71:60] = in_4[71:60] / Quant[4][5];
		if(in_4[59:48] > 12'b011111111111)
		begin
			q_4[59:48] = ((in_4[59:48]^12'b111111111111)+1) / Quant[4][4];
			if (q_4[59:48] >0) q_4[59:48] =(q_4[59:48]^12'b111111111111)+1;
		end
		else q_4[59:48] = in_4[59:48] / Quant[4][4];
		if(in_4[47:36] > 12'b011111111111)
		begin
			q_4[47:36] = ((in_4[47:36]^12'b111111111111)+1) / Quant[4][3];
			if (q_4[47:36] >0) q_4[47:36] =(q_4[47:36]^12'b111111111111)+1;
		end
		else q_4[47:36] = in_4[47:36] / Quant[4][3];
		if(in_4[35:24] > 12'b011111111111)
		begin
			q_4[35:24] = ((in_4[35:24]^12'b111111111111)+1) / Quant[4][2];
			if (q_4[35:24] >0) q_4[35:24] =(q_4[35:24]^12'b111111111111)+1;
		end
		else q_4[35:24] = in_4[35:24] / Quant[4][2];
		if(in_4[23:12] > 12'b011111111111)
		begin
			q_4[23:12] = ((in_4[23:12]^12'b111111111111)+1) / Quant[4][1];
			if (q_4[23:12] >0) q_4[23:12] =(q_4[23:12]^12'b111111111111)+1;
		end
		else q_4[23:12] = in_4[23:12] / Quant[4][1];
		if(in_4[11:0]  > 12'b011111111111)
		begin
			q_4[11:0]  = ((in_4[11:0] ^12'b111111111111)+1) / Quant[4][0];
			if (q_4[11:0]  >0) q_4[11:0]  =(q_4[11:0] ^12'b111111111111)+1;
		end
		else q_4[11:0]  = in_4[11:0]  / Quant[4][0];
		
		if(in_5[95:84] > 12'b011111111111)
		begin
			q_5[95:84] = ((in_5[95:84]^12'b111111111111)+1) / Quant[5][7];
			if (q_5[95:84] >0) q_5[95:84] =(q_5[95:84]^12'b111111111111)+1;
		end
		else q_5[95:84] = in_5[95:84] / Quant[5][7];
		if(in_5[83:72] > 12'b011111111111)
		begin
			q_5[83:72] = ((in_5[83:72]^12'b111111111111)+1) / Quant[5][6];
			if (q_5[83:72] >0) q_5[83:72] =(q_5[83:72]^12'b111111111111)+1;
		end
		else q_5[83:72] = in_5[83:72] / Quant[5][6];
		if(in_5[71:60] > 12'b011111111111)
		begin
			q_5[71:60] = ((in_5[71:60]^12'b111111111111)+1) / Quant[5][5];
			if (q_5[71:60] >0) q_5[71:60] =(q_5[71:60]^12'b111111111111)+1;
		end
		else q_5[71:60] = in_5[71:60] / Quant[5][5];
		if(in_5[59:48] > 12'b011111111111)
		begin
			q_5[59:48] = ((in_5[59:48]^12'b111111111111)+1) / Quant[5][4];
			if (q_5[59:48] >0) q_5[59:48] =(q_5[59:48]^12'b111111111111)+1;
		end
		else q_5[59:48] = in_5[59:48] / Quant[5][4];
		if(in_5[47:36] > 12'b011111111111)
		begin
			q_5[47:36] = ((in_5[47:36]^12'b111111111111)+1) / Quant[5][3];
			if (q_5[47:36] >0) q_5[47:36] =(q_5[47:36]^12'b111111111111)+1;
		end
		else q_5[47:36] = in_5[47:36] / Quant[5][3];
		if(in_5[35:24] > 12'b011111111111)
		begin
			q_5[35:24] = ((in_5[35:24]^12'b111111111111)+1) / Quant[5][2];
			if (q_5[35:24] >0) q_5[35:24] =(q_5[35:24]^12'b111111111111)+1;
		end
		else q_5[35:24] = in_5[35:24] / Quant[5][2];
		if(in_5[23:12] > 12'b011111111111)
		begin
			q_5[23:12] = ((in_5[23:12]^12'b111111111111)+1) / Quant[5][1];
			if (q_5[23:12] >0) q_5[23:12] =(q_5[23:12]^12'b111111111111)+1;
		end
		else q_5[23:12] = in_5[23:12] / Quant[5][1];
		if(in_5[11:0]  > 12'b011111111111)
		begin
			q_5[11:0]  = ((in_5[11:0] ^12'b111111111111)+1) / Quant[5][0];
			if (q_5[11:0]  >0) q_5[11:0]  =(q_5[11:0] ^12'b111111111111)+1;
		end
		else q_5[11:0]  = in_5[11:0]  / Quant[5][0];
		
		if(in_6[95:84] > 12'b011111111111)
		begin
			q_6[95:84] = ((in_6[95:84]^12'b111111111111)+1) / Quant[6][7];
			if (q_6[95:84] >0) q_6[95:84] =(q_6[95:84]^12'b111111111111)+1;
		end
		else q_6[95:84] = in_6[95:84] / Quant[6][7];
		if(in_6[83:72] > 12'b011111111111)
		begin
			q_6[83:72] = ((in_6[83:72]^12'b111111111111)+1) / Quant[6][6];
			if (q_6[83:72] >0) q_6[83:72] =(q_6[83:72]^12'b111111111111)+1;
		end
		else q_6[83:72] = in_6[83:72] / Quant[6][6];
		if(in_6[71:60] > 12'b011111111111)
		begin
			q_6[71:60] = ((in_6[71:60]^12'b111111111111)+1) / Quant[6][5];
			if (q_6[71:60] >0) q_6[71:60] =(q_6[71:60]^12'b111111111111)+1;
		end
		else q_6[71:60] = in_6[71:60] / Quant[6][5];
		if(in_6[59:48] > 12'b011111111111)
		begin
			q_6[59:48] = ((in_6[59:48]^12'b111111111111)+1) / Quant[6][4];
			if (q_6[59:48] >0) q_6[59:48] =(q_6[59:48]^12'b111111111111)+1;
		end
		else q_6[59:48] = in_6[59:48] / Quant[6][4];
		if(in_6[47:36] > 12'b011111111111)
		begin
			q_6[47:36] = ((in_6[47:36]^12'b111111111111)+1) / Quant[6][3];
			if (q_6[47:36] >0) q_6[47:36] =(q_6[47:36]^12'b111111111111)+1;
		end
		else q_6[47:36] = in_6[47:36] / Quant[6][3];
		if(in_6[35:24] > 12'b011111111111)
		begin
			q_6[35:24] = ((in_6[35:24]^12'b111111111111)+1) / Quant[6][2];
			if (q_6[35:24] >0) q_6[35:24] =(q_6[35:24]^12'b111111111111)+1;
		end
		else q_6[35:24] = in_6[35:24] / Quant[6][2];
		if(in_6[23:12] > 12'b011111111111)
		begin
			q_6[23:12] = ((in_6[23:12]^12'b111111111111)+1) / Quant[6][1];
			if (q_6[23:12] >0) q_6[23:12] =(q_6[23:12]^12'b111111111111)+1;
		end
		else q_6[23:12] = in_6[23:12] / Quant[6][1];
		if(in_6[11:0]  > 12'b011111111111)
		begin
			q_6[11:0]  = ((in_6[11:0] ^12'b111111111111)+1) / Quant[6][0];
			if (q_6[11:0]  >0) q_6[11:0]  =(q_6[11:0] ^12'b111111111111)+1;
		end
		else q_6[11:0]  = in_6[11:0]  / Quant[6][0];
		
		if(in_7[95:84] > 12'b011111111111)
		begin
			q_7[95:84] = ((in_7[95:84]^12'b111111111111)+1) / Quant[7][7];
			if (q_7[95:84] >0) q_7[95:84] =(q_7[95:84]^12'b111111111111)+1;
		end
		else q_7[95:84] = in_7[95:84] / Quant[7][7];
		if(in_7[83:72] > 12'b011111111111)
		begin
			q_7[83:72] = ((in_7[83:72]^12'b111111111111)+1) / Quant[7][6];
			if (q_7[83:72] >0) q_7[83:72] =(q_7[83:72]^12'b111111111111)+1;
		end
		else q_7[83:72] = in_7[83:72] / Quant[7][6];
		if(in_7[71:60] > 12'b011111111111)
		begin
			q_7[71:60] = ((in_7[71:60]^12'b111111111111)+1) / Quant[7][5];
			if (q_7[71:60] >0) q_7[71:60] =(q_7[71:60]^12'b111111111111)+1;
		end
		else q_7[71:60] = in_7[71:60] / Quant[7][5];
		if(in_7[59:48] > 12'b011111111111)
		begin
			q_7[59:48] = ((in_7[59:48]^12'b111111111111)+1) / Quant[7][4];
			if (q_7[59:48] >0) q_7[59:48] =(q_7[59:48]^12'b111111111111)+1;
		end
		else q_7[59:48] = in_7[59:48] / Quant[7][4];
		if(in_7[47:36] > 12'b011111111111)
		begin
			q_7[47:36] = ((in_7[47:36]^12'b111111111111)+1) / Quant[7][3];
			if (q_7[47:36] >0) q_7[47:36] =(q_7[47:36]^12'b111111111111)+1;
		end
		else q_7[47:36] = in_7[47:36] / Quant[7][3];
		if(in_7[35:24] > 12'b011111111111)
		begin
			q_7[35:24] = ((in_7[35:24]^12'b111111111111)+1) / Quant[7][2];
			if (q_7[35:24] >0) q_7[35:24] =(q_7[35:24]^12'b111111111111)+1;
		end
		else q_7[35:24] = in_7[35:24] / Quant[7][2];
		if(in_7[23:12] > 12'b011111111111)
		begin
			q_7[23:12] = ((in_7[23:12]^12'b111111111111)+1) / Quant[7][1];
			if (q_7[23:12] >0) q_7[23:12] =(q_7[23:12]^12'b111111111111)+1;
		end
		else q_7[23:12] = in_7[23:12] / Quant[7][1];
		if(in_7[11:0]  > 12'b011111111111)
		begin
			q_7[11:0]  = ((in_7[11:0] ^12'b111111111111)+1) / Quant[7][0];
			if (q_7[11:0]  >0) q_7[11:0]  =(q_7[11:0] ^12'b111111111111)+1;
		end
		else q_7[11:0]  = in_7[11:0]  / Quant[7][0];
	end
endmodule
