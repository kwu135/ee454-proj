`timescale 1 ns / 100 ps

module tb_generateDCT();

reg[63:0] pixels_0;
reg[63:0] pixels_1;
reg[63:0] pixels_2;
reg[63:0] pixels_3;
reg[63:0] pixels_4;
reg[63:0] pixels_5;
reg[63:0] pixels_6;
reg[63:0] pixels_7;

reg Clk;
reg Reset;
wire[95:0] dct_0;
wire[95:0] dct_1;
wire[95:0] dct_2;
wire[95:0] dct_3;
wire[95:0] dct_4;
wire[95:0] dct_5;
wire[95:0] dct_6;
wire[95:0] dct_7;

wire Done;
parameter CLK_PERIOD=2;
always 	#(CLK_PERIOD/2) Clk=~Clk;

initial 
begin
Clk=0;
Reset =0;

pixels_0 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_1 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_2 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_3 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_4 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_5 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_6 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

pixels_7 = 
8'b000000000000 << 56 |
8'b000000000000 << 48 |
8'b000000000000 << 40 |
8'b000000000000 << 32 |
8'b000000000000 << 24 |
8'b000000000000 << 16 |
8'b000000000000 << 8 |
8'b000000000000;

#(CLK_PERIOD)
Reset = 1;
#(CLK_PERIOD)
Reset = 0;
#(CLK_PERIOD * 400)
$stop;
end

generateDCT dct(pixels_0, pixels_1, pixels_2, pixels_3, pixels_4,
	pixels_5, pixels_6, pixels_7, Clk, Reset, dct_0, dct_1, dct_2, dct_3,
	dct_4, dct_5, dct_6, dct_7, Done);
endmodule